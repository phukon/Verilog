//-----------------------------------------------------------------------------
//
// Title       : multiplier
// Design      : gates
// Author      : 
// Company     : 
//
//-----------------------------------------------------------------------------
//
// File        : d:\desktop files\core 2 (exim)\Projects\Aldec\Diversity_techniques\gates\src\multiplier.v
// Generated   : Wed Aug 31 14:39:09 2022
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {multiplier}}
module multiplier ( y1 ,y2 ,out );

input wire y1, y2 ;

output out ;
assign out = y1 * y2;  
wire out ;
//}} End of automatically maintained section

// -- Enter your statements here -- //

endmodule
